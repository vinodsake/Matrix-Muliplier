/**********************************************************************
* File Name	: package.sv
* Description 	: Includes common variables, parameters, tasks/funcs
* Creation Date : 06-12-2020
* Last Modified : Sun 17 Jan 2021 04:48:08 PM PST
* Author 	: Vinod Sake
* Email 	: vinodsake042@gmail.com
* GitHub	: github.com/vinodsake
**********************************************************************/
`ifndef PACKAGE_DONE
`define PACKAGE_DONE
package project_pkg;
	parameter MSB = 32;
endpackage : project_pkg
`endif
